ampli
i1 0 1 ac 1
r1 1 0 820000
r2 2 1 100
r3 2 0 10400
c1 2 0 57e-12
c2 2 3 4.5e-12
g1 3 0 2 0 0.038
r4 3 0 4700
r5 3 0 820k
.ac dec 1000 1k 10Meg
.probe
.end

